`define IDLE   3'b000
`define START  3'b001 
`define DATA   3'b011
`define PARITY 3'b010
`define STOP   3'b110